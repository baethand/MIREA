library verilog;
use verilog.vl_types.all;
entity Q41_vlg_vec_tst is
end Q41_vlg_vec_tst;
