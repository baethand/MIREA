library verilog;
use verilog.vl_types.all;
entity Q42_vlg_vec_tst is
end Q42_vlg_vec_tst;
